----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:04:21 10/24/2022 
-- Design Name: 
-- Module Name:    Product_Register - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Product_Register is

generic (n: integer := 16);

port(
	clk, pload : in std_logic;
	D_in       : in std_logic_vector(n-1 downto 0);
	Q_out      : out std_logic_vector(n-1 downto 0) 
	

);
end Product_Register;

architecture Behavioral of Product_Register is

begin

register_proc: process (clk)
	begin
	 
	 if (rising_edge(clk)) then
	   if (pload = '1') then
		   Q_out <= D_in;
		end if;	
	 end if;
end process;
	 

end Behavioral;

